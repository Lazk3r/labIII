library verilog;
use verilog.vl_types.all;
entity MOORE_TEST1_vlg_vec_tst is
end MOORE_TEST1_vlg_vec_tst;
