-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Jun 21 11:08:08 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mealy IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        X : IN STD_LOGIC := '0';
        Z : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END mealy;

ARCHITECTURE BEHAVIOR OF mealy IS
    TYPE type_fstate IS (state0,state1,state2,state3,state4,state5,state6,state7,state8,state9,state10);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,X)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state0;
            Z <= "00";
        ELSE
            Z <= "00";
            CASE fstate IS
                WHEN state0 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state0;
                    END IF;

                    Z <= "00";
                WHEN state1 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    Z <= "00";
                WHEN state2 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    Z <= "00";
                WHEN state3 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    IF ((X = '0')) THEN
                        Z <= "00";
                    ELSIF ((X = '1')) THEN
                        Z <= "10";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= "00";
                    END IF;
                WHEN state4 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state8;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    IF ((X = '0')) THEN
                        Z <= "01";
                    ELSIF ((X = '1')) THEN
                        Z <= "00";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= "00";
                    END IF;
                WHEN state5 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    Z <= "00";
                WHEN state6 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    Z <= "00";
                WHEN state7 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state8;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    IF ((X = '1')) THEN
                        Z <= "00";
                    ELSIF ((X = '0')) THEN
                        Z <= "01";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= "00";
                    END IF;
                WHEN state8 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state8;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    Z <= "01";
                WHEN state9 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state8;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    Z <= "01";
                WHEN state10 =>
                    IF ((X = '0')) THEN
                        reg_fstate <= state1;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    IF ((X = '1')) THEN
                        Z <= "10";
                    ELSIF ((X = '0')) THEN
                        Z <= "00";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= "00";
                    END IF;
                WHEN OTHERS => 
                    Z <= "XX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
